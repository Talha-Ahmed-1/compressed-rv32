module CompressedDecoder(
  input         clock,
  input         reset,
  input  [31:0] io_instIn,
  output [31:0] io_instOut,
  output        io_compressed
);
  wire [3:0] _GEN_0 = {{1'd0}, io_instIn[4:2]}; // @[CompressedDecoder.scala 51:27]
  wire [3:0] _RS1_T_2 = _GEN_0 + 4'h8; // @[CompressedDecoder.scala 51:27]
  wire [3:0] _GEN_1 = {{1'd0}, io_instIn[9:7]}; // @[CompressedDecoder.scala 53:30]
  wire [3:0] _RD_RS2_T_2 = _GEN_1 + 4'h8; // @[CompressedDecoder.scala 53:30]
  wire [15:0] _T_1 = io_instIn[15:0] & 16'he003; // @[CompressedDecoder.scala 66:26]
  wire  _T_2 = 16'h4000 == _T_1; // @[CompressedDecoder.scala 66:26]
  wire  hi_hi_hi = io_instIn[5]; // @[CompressedDecoder.scala 55:32]
  wire [2:0] hi_hi_lo = io_instIn[12:10]; // @[CompressedDecoder.scala 55:46]
  wire  hi_lo_hi = io_instIn[6]; // @[CompressedDecoder.scala 55:64]
  wire [4:0] RS1 = {{1'd0}, _RS1_T_2}; // @[CompressedDecoder.scala 50:19 CompressedDecoder.scala 51:9]
  wire [4:0] RD_RS2 = {{1'd0}, _RD_RS2_T_2}; // @[CompressedDecoder.scala 52:22 CompressedDecoder.scala 53:12]
  wire [19:0] _T_3 = {hi_hi_hi,hi_hi_lo,hi_lo_hi,1'h0,RD_RS2,2'h2,RS1,2'h3}; // @[Cat.scala 30:58]
  wire  _T_6 = 16'hc000 == _T_1; // @[CompressedDecoder.scala 70:26]
  wire  hi_hi_lo_1 = io_instIn[12]; // @[CompressedDecoder.scala 56:58]
  wire [1:0] lo_hi_hi_lo = io_instIn[11:10]; // @[CompressedDecoder.scala 56:96]
  wire [24:0] _T_7 = {1'h0,hi_hi_hi,hi_hi_lo_1,RS1,RD_RS2,2'h2,lo_hi_hi_lo,hi_lo_hi,7'h23}; // @[Cat.scala 30:58]
  wire [15:0] _T_9 = io_instIn[15:0] & 16'hfc63; // @[CompressedDecoder.scala 91:26]
  wire  _T_10 = 16'h8c61 == _T_9; // @[CompressedDecoder.scala 91:26]
  wire [25:0] _T_11 = {1'h0,RD_RS2,RS1,3'h7,RD_RS2,7'h33}; // @[Cat.scala 30:58]
  wire  _T_14 = 16'h8c41 == _T_9; // @[CompressedDecoder.scala 92:26]
  wire [25:0] _T_15 = {1'h0,RD_RS2,RS1,3'h6,RD_RS2,7'h33}; // @[Cat.scala 30:58]
  wire  _T_18 = 16'h8c21 == _T_9; // @[CompressedDecoder.scala 93:26]
  wire [25:0] _T_19 = {1'h0,RD_RS2,RS1,3'h4,RD_RS2,7'h33}; // @[Cat.scala 30:58]
  wire  _T_22 = 16'h8c01 == _T_9; // @[CompressedDecoder.scala 94:26]
  wire [30:0] _T_23 = {6'h20,RD_RS2,RS1,3'h0,RD_RS2,7'h33}; // @[Cat.scala 30:58]
  wire  _T_26 = 16'h1 == io_instIn[15:0]; // @[CompressedDecoder.scala 95:26]
  wire  _T_29 = 16'h9002 == io_instIn[15:0]; // @[CompressedDecoder.scala 96:26]
  wire  _T_32 = 16'h0 == io_instIn[15:0]; // @[CompressedDecoder.scala 97:26]
  wire [31:0] _io_instOut_T = _T_32 ? 32'h0 : io_instIn; // @[Mux.scala 98:16]
  wire [31:0] _io_instOut_T_1 = _T_29 ? 32'h100073 : _io_instOut_T; // @[Mux.scala 98:16]
  wire [31:0] _io_instOut_T_2 = _T_26 ? 32'h13 : _io_instOut_T_1; // @[Mux.scala 98:16]
  wire [31:0] _io_instOut_T_3 = _T_22 ? {{1'd0}, _T_23} : _io_instOut_T_2; // @[Mux.scala 98:16]
  wire [31:0] _io_instOut_T_4 = _T_18 ? {{6'd0}, _T_19} : _io_instOut_T_3; // @[Mux.scala 98:16]
  wire [31:0] _io_instOut_T_5 = _T_14 ? {{6'd0}, _T_15} : _io_instOut_T_4; // @[Mux.scala 98:16]
  wire [31:0] _io_instOut_T_6 = _T_10 ? {{6'd0}, _T_11} : _io_instOut_T_5; // @[Mux.scala 98:16]
  wire [31:0] _io_instOut_T_7 = _T_6 ? {{7'd0}, _T_7} : _io_instOut_T_6; // @[Mux.scala 98:16]
  assign io_instOut = _T_2 ? {{12'd0}, _T_3} : _io_instOut_T_7; // @[Mux.scala 98:16]
  assign io_compressed = io_instIn != io_instOut; // @[CompressedDecoder.scala 100:32]
endmodule
